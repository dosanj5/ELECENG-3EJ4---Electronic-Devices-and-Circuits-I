** Profile: "SCHEMATIC1-step1_3"  [ c:\users\dosanj5\onedrive - mcmaster university\school files\2025 - 2026\elec 3ej4\lab 4\pspice\3ej4 lab 4-PSpiceFiles\SCHEMATIC1\step1_3.sim ] 

** Creating circuit file "step1_3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\dosanj5\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "C:\Users\dosanj5\OneDrive - McMaster University\School Files\2025 - 2026\ELEC 3EJ4\Model Parts\My2N3906.LIB" 
.lib "C:\Users\dosanj5\OneDrive - McMaster University\School Files\2025 - 2026\ELEC 3EJ4\Model Parts\My2N3904.LIB" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 101 100Hz 100kHz
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
