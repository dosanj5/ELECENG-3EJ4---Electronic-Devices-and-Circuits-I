** Profile: "PART3-dc_sweep_pt3"  [ C:\Users\dosanj5\OneDrive - McMaster University\School Files\2025 - 2026\ELEC 3EJ4\Lab 1\PSpice\3EJ4 Lab 1-PSpiceFiles\PART3\dc_sweep_pt3.sim ] 

** Creating circuit file "dc_sweep_pt3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\dosanj5\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "C:\Users\dosanj5\OneDrive - McMaster University\School Files\2025 - 2026\ELEC 3EJ4\Model Parts\My2N3906.LIB" 
.lib "C:\Users\dosanj5\OneDrive - McMaster University\School Files\2025 - 2026\ELEC 3EJ4\Model Parts\My2N3904.LIB" 
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VCC -5 5 0.05 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\PART3.net" 


.END
